library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Memoria is
	 generic(
			f_reloj: integer:= 12000000;
			f_media_onda:integer:= 308; 
			bits_salida: integer:= 12;
			direcciones: integer:= 500);
    Port ( 
			  Clk : in  STD_LOGIC;
           SALIDA : out  STD_LOGIC_VECTOR (bits_salida-1 downto 0));
			  
end Memoria;

architecture Behavioral of Memoria is

	 type rom_type is array (direcciones-1 downto 0) of std_logic_vector (bits_salida-1 downto 0);                 
    constant ROM : rom_type:= (
"100000000000","111111111111","111111111111","111111111111","111111111111","111111111110","111111111110","111111111110","111111111101","111111111100",
"111111111011","111111111011","111111111010","111111111001","111111111000","111111110110","111111110101","111111110100","111111110010","111111110001",
"111111101111","111111101110","111111101100","111111101010","111111101000","111111100110","111111100100","111111100010","111111100000","111111011101",
"111111011011","111111011001","111111010110","111111010011","111111010001","111111001110","111111001011","111111001000","111111000101","111111000010",
"111110111111","111110111100","111110111000","111110110101","111110110001","111110101110","111110101010","111110100110","111110100011","111110011111",
"111110011011","111110010111","111110010011","111110001111","111110001010","111110000110","111110000010","111101111101","111101111000","111101110100",
"111101101111","111101101010","111101100101","111101100001","111101011011","111101010110","111101010001","111101001100","111101000111","111101000001",
"111100111100","111100110110","111100110001","111100101011","111100100101","111100011111","111100011010","111100010100","111100001101","111100000111",
"111100000001","111011111011","111011110101","111011101110","111011101000","111011100001","111011011011","111011010100","111011001101","111011000110",
"111010111111","111010111000","111010110001","111010101010","111010100011","111010011100","111010010101","111010001101","111010000110","111001111110",
"111001110111","111001101111","111001101000","111001100000","111001011000","111001010000","111001001000","111001000000","111000111000","111000110000",
"111000101000","111000011111","111000010111","111000001111","111000000110","110111111110","110111110101","110111101101","110111100100","110111011011",
"110111010010","110111001001","110111000001","110110111000","110110101110","110110100101","110110011100","110110010011","110110001010","110110000000",
"110101110111","110101101110","110101100100","110101011011","110101010001","110101000111","110100111110","110100110100","110100101010","110100100000",
"110100010110","110100001100","110100000010","110011111000","110011101110","110011100100","110011011010","110011001111","110011000101","110010111011",
"110010110000","110010100110","110010011011","110010010001","110010000110","110001111011","110001110001","110001100110","110001011011","110001010000",
"110001000101","110000111010","110000110000","110000100100","110000011001","110000001110","110000000011","101111111000","101111101101","101111100010",
"101111010110","101111001011","101111000000","101110110100","101110101001","101110011101","101110010010","101110000110","101101111011","101101101111",
"101101100011","101101011000","101101001100","101101000000","101100110100","101100101000","101100011101","101100010001","101100000101","101011111001",
"101011101101","101011100001","101011010101","101011001001","101010111101","101010110001","101010100100","101010011000","101010001100","101010000000",
"101001110011","101001100111","101001011011","101001001111","101001000010","101000110110","101000101001","101000011101","101000010001","101000000100",
"100111111000","100111101011","100111011111","100111010010","100111000101","100110111001","100110101100","100110100000","100110010011","100110000110",
"100101111010","100101101101","100101100000","100101010100","100101000111","100100111010","100100101101","100100100001","100100010100","100100000111",
"100011111010","100011101101","100011100001","100011010100","100011000111","100010111010","100010101101","100010100001","100010010100","100010000111",
"100001111010","100001101101","100001100000","100001010011","100001000110","100000111010","100000101101","100000100000","100000010011","100000000110",
"011111111001","011111101100","011111011111","011111010010","011111000101","011110111001","011110101100","011110011111","011110010010","011110000101",
"011101111000","011101101011","011101011110","011101010010","011101000101","011100111000","011100101011","011100011110","011100010010","011100000101",
"011011111000","011011101011","011011011110","011011010010","011011000101","011010111000","011010101011","011010011111","011010010010","011010000101",
"011001111001","011001101100","011001011111","011001010011","011001000110","011000111010","011000101101","011000100000","011000010100","011000000111",
"010111111011","010111101110","010111100010","010111010110","010111001001","010110111101","010110110000","010110100100","010110011000","010110001100",
"010101111111","010101110011","010101100111","010101011011","010101001110","010101000010","010100110110","010100101010","010100011110","010100010010",
"010100000110","010011111010","010011101110","010011100010","010011010111","010011001011","010010111111","010010110011","010010100111","010010011100",
"010010010000","010010000100","010001111001","010001101101","010001100010","010001010110","010001001011","010000111111","010000110100","010000101001",
"010000011101","010000010010","010000000111","001111111100","001111110001","001111100110","001111011011","001111001111","001111000101","001110111010",
"001110101111","001110100100","001110011001","001110001110","001110000100","001101111001","001101101110","001101100100","001101011001","001101001111",
"001101000100","001100111010","001100110000","001100100101","001100011011","001100010001","001100000111","001011111101","001011110011","001011101001",
"001011011111","001011010101","001011001011","001011000001","001010111000","001010101110","001010100100","001010011011","001010010001","001010001000",
"001001111111","001001110101","001001101100","001001100011","001001011010","001001010001","001001000111","001000111110","001000110110","001000101101",
"001000100100","001000011011","001000010010","001000001010","001000000001","000111111001","000111110000","000111101000","000111100000","000111010111",
"000111001111","000111000111","000110111111","000110110111","000110101111","000110100111","000110011111","000110010111","000110010000","000110001000",
"000110000001","000101111001","000101110010","000101101010","000101100011","000101011100","000101010101","000101001110","000101000111","000101000000",
"000100111001","000100110010","000100101011","000100100100","000100011110","000100010111","000100010001","000100001010","000100000100","000011111110",
"000011111000","000011110010","000011101011","000011100101","000011100000","000011011010","000011010100","000011001110","000011001001","000011000011",
"000010111110","000010111000","000010110011","000010101110","000010101001","000010100100","000010011110","000010011010","000010010101","000010010000",
"000010001011","000010000111","000010000010","000001111101","000001111001","000001110101","000001110000","000001101100","000001101000","000001100100",
"000001100000","000001011100","000001011001","000001010101","000001010001","000001001110","000001001010","000001000111","000001000011","000001000000",
"000000111101","000000111010","000000110111","000000110100","000000110001","000000101110","000000101100","000000101001","000000100110","000000100100",
"000000100010","000000011111","000000011101","000000011011","000000011001","000000010111","000000010101","000000010011","000000010001","000000010000",
"000000001110","000000001101","000000001011","000000001010","000000001001","000000000111","000000000110","000000000101","000000000100","000000000100",
"000000000011","000000000010","000000000001","000000000001","000000000001","000000000000","000000000000","000000000000","000000000000","000000000000"
	  );
	 
	 signal contador: integer range 0 to f_media_onda:= 0;
	 signal dir: integer range 0 to direcciones-1:= 0;
	 signal hight_low: std_logic:= '0';
	 signal cambio: std_logic:= '0';
	 
begin

	control: process(CLK)
	begin
		if (rising_edge(CLK)) then
			if (contador < f_media_onda) then
				contador <= contador + 1;
			else
				contador <= 0;
				cambio <= not cambio;
				if (hight_low = '0') then 
					if (dir < direcciones-1) then 
						dir <= dir + 1;
					else
						hight_low <= '1';
					end if;
				elsif (hight_low = '1') then 
					if (dir > 0) then 
						dir <= dir - 1;
					else
						hight_low <= '0';
					end if;
				end if;
			end if;
		end if;
	end process control;
	
	parpadeo: process(cambio,dir)
	begin
		SALIDA <= ROM(dir);
	end process parpadeo;
	
end Behavioral;

